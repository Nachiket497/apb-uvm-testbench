package enums;

  typedef enum {
    IDLE,
    SETUP,
    ACCESS
  } apb_state;

endpackage

